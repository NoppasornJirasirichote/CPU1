`timescale 1ns / 1ps

module OR(
    input A,
	 input B,
	 output out);
	 
	 or(out,A,B);
	 
endmodule

`timescale 1ns / 1ps

module AND(
    input A,
	 input B,
	 output out);
	 
	 and(out,A,B);


endmodule

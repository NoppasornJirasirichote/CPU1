`timescale 1ns / 1ps

module sub(
    input [7:0]A,
	 input [7:0]B,
	 output [7:0]out);
	 
	 assign out = A-B;


endmodule

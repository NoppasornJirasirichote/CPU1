`timescale 1ns / 1ps

module Main(
    );


endmodule
